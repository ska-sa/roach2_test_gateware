module qdrc_infrastructure(
    /* general signals */
    clk0,
    clk180,
    clk270,
    /* external signals */
    qdr_d,
    qdr_q,
    qdr_sa,
    qdr_w_n,
    qdr_r_n,
    qdr_dll_off_n,
    qdr_k,
    qdr_k_n,
    /* phy->external signals */
    qdr_d_rise,
    qdr_d_fall,
    qdr_q_rise,
    qdr_q_fall,
    qdr_sa_buf,
    qdr_w_n_buf,
    qdr_r_n_buf,
    qdr_dll_off_n_buf,
    /* phy training signals */
    dly_clk,
    dly_inc_dec_n,
    dly_en,
    dly_rst       
  );
  parameter DATA_WIDTH     = 36;
  parameter ADDR_WIDTH     = 21;
  parameter CLK_FREQ       = 200;

  input clk0,   clk180,   clk270;

  output [DATA_WIDTH - 1:0] qdr_d;
  input  [DATA_WIDTH - 1:0] qdr_q;
  output [ADDR_WIDTH - 1:0] qdr_sa;
  output qdr_w_n;
  output qdr_r_n;
  output qdr_dll_off_n;
  output qdr_k, qdr_k_n;
  
  input  [DATA_WIDTH - 1:0] qdr_d_rise;
  input  [DATA_WIDTH - 1:0] qdr_d_fall;
  output [DATA_WIDTH - 1:0] qdr_q_rise;
  output [DATA_WIDTH - 1:0] qdr_q_fall;
  input  [ADDR_WIDTH - 1:0] qdr_sa_buf;
  input  qdr_w_n_buf, qdr_r_n_buf;
  input  qdr_dll_off_n_buf;

  input  dly_clk;
  input  [DATA_WIDTH - 1:0] dly_inc_dec_n;
  input  [DATA_WIDTH - 1:0] dly_en;
  input  [DATA_WIDTH - 1:0] dly_rst;       

  /******************* QDR_K and QDR_K_N ********************
   * The clock is generated by an ODDR. This is done
   * to so the latency introduced by the ODDR on the data
   * line is introduced into the clock generation.
   * The clock uses clk0 while all other signals use clk270.
   */

  ODDR #(
    .DDR_CLK_EDGE ("SAME_EDGE"),
    .INIT         (1'b1),
    .SRTYPE       ("SYNC")
  ) ODDR_qdr_k (
    .Q  (qdr_k),
    .C  (clk0),
    .CE (1'b1),
    .D1 (1'b1), //Rising Edge
    .D2 (1'b0), //Falling Edge
    .R  (1'b0),
    .S  (1'b0)
  );

  /* same as qdr_k -> just inverted */
  ODDR #(
    .DDR_CLK_EDGE ("SAME_EDGE"),
    .INIT         (1'b1),
    .SRTYPE       ("SYNC")
  ) ODDR_qdr_k_n (
    .Q  (qdr_k_n),
    .C  (clk0),
    .CE (1'b1),
    .D1 (1'b0), //Rising Edge
    .D2 (1'b1), //Falling Edge
    .R  (1'b0),
    .S  (1'b0)
  );

  /******************* SDR Control Signals ********************
   *
   */

  reg [ADDR_WIDTH - 1:0] qdr_sa_reg;
  reg qdr_w_n_reg;
  reg qdr_r_n_reg;

  /* This signals are all sliced so use the register in the slice */

  always @(posedge clk0) begin 
    qdr_sa_reg        <= qdr_sa_buf;
    qdr_w_n_reg       <= qdr_w_n_buf;
    qdr_r_n_reg       <= qdr_r_n_buf;
  end

  reg [ADDR_WIDTH - 1:0] qdr_sa_reg0;
  reg qdr_w_n_reg0;
  reg qdr_r_n_reg0;

  always @(posedge clk180) begin 
  /* Add delay to ease timing */
    qdr_sa_reg0        <= qdr_sa_reg;
    qdr_w_n_reg0       <= qdr_w_n_reg;
    qdr_r_n_reg0       <= qdr_r_n_reg;
  end

  reg [ADDR_WIDTH - 1:0] qdr_sa_iob;
  reg qdr_w_n_iob;
  reg qdr_r_n_iob;
  //synthesis attribute IOB of qdr_sa_iob        is "TRUE"
  //synthesis attribute IOB of qdr_w_n_iob       is "TRUE"
  //synthesis attribute IOB of qdr_r_n_iob       is "TRUE"


  always @(posedge clk180) begin 
  /* Add delay to ease timing */
    qdr_sa_iob        <= qdr_sa_reg0;
    qdr_w_n_iob       <= qdr_w_n_reg0;
    qdr_r_n_iob       <= qdr_r_n_reg0;
  end

  OBUF OBUF_addr[ADDR_WIDTH - 1:0](
    .I (qdr_sa_iob),
    .O (qdr_sa)
  );

  OBUF OBUF_w_n(
    .I (qdr_w_n_iob),
    .O (qdr_w_n)
  );

  OBUF OBUF_r_n(
    .I (qdr_r_n_iob),
    .O (qdr_r_n)
  );

  OBUF OBUF_dll_off_n(
    .I (qdr_dll_off_n_buf),
    .O (qdr_dll_off_n)
  );


  /******************* DDR Data Outputs ********************
   *
   */

  reg [DATA_WIDTH - 1:0] qdr_d_rise_reg0;
  reg [DATA_WIDTH - 1:0] qdr_d_fall_reg0;

  always @(posedge clk0) begin
  /* Delay the write data by one cycle (qdr protocol,
   * requires datat to lag control*/
    qdr_d_rise_reg0     <= qdr_d_rise;
    qdr_d_fall_reg0     <= qdr_d_fall;
  end

  reg [DATA_WIDTH - 1:0] qdr_d_rise_reg1;
  reg [DATA_WIDTH - 1:0] qdr_d_fall_reg1;

  always @(posedge clk0) begin
  /* Delay to match the extra cycle on control lines 
   * due to extra iob delay route*/
    qdr_d_rise_reg1     <= qdr_d_rise_reg0;
    qdr_d_fall_reg1     <= qdr_d_fall_reg0;
  end


  reg [DATA_WIDTH - 1:0] qdr_d_rise_reg;
  reg [DATA_WIDTH - 1:0] qdr_d_fall_reg;

  always @(posedge clk270) begin
  /* Sample DDR signals onto clk270 domain.
   * The 270 clock is used to let the data lead the clock by
   * 90 degrees behind the clock. The signals are registered
   * to ease timing requirements.
   */
    qdr_d_rise_reg     <= qdr_d_rise_reg1;
    qdr_d_fall_reg     <= qdr_d_fall_reg1;
  end

  ODDR #(
    .DDR_CLK_EDGE ("SAME_EDGE"),
    .INIT         (1'b1),
    .SRTYPE       ("SYNC")
  ) ODDR_qdr_d [DATA_WIDTH - 1:0] (
    .Q  (qdr_d),
    .C  (clk270),
    .CE (1'b1),
    .D1 (qdr_d_rise_reg), //Rising Edge
    .D2 (qdr_d_fall_reg), //Falling Edge
    .R  (1'b0),
    .S  (1'b0)
  );

  /******************* DDR Data Inputs ********************
   * IODELAY for training
   */
 
  wire [DATA_WIDTH - 1:0] qdr_q_ibuf;
  wire [DATA_WIDTH - 1:0] qdr_q_iodelay;

  IBUF ibuf_qdrq [DATA_WIDTH - 1:0](
    .I (qdr_q),
    .O (qdr_q_ibuf)
  );

  IODELAY #(
    .DELAY_SRC        ("I"),
    .IDELAY_TYPE      ("VARIABLE"),
    .REFCLK_FREQUENCY (200.0)
  ) IODELAY_qdrq [DATA_WIDTH - 1:0] (
    .C       (dly_clk),
    .CE      (dly_en),
    .DATAIN  (1'b0),
    .IDATAIN (qdr_q_ibuf),
    .INC     (dly_inc_dec_n),
    .ODATAIN (),
    .RST     (dly_rst),
    .T       (1'b0),
    .DATAOUT (qdr_q_iodelay)
  );

  wire [DATA_WIDTH - 1:0] qdr_q_rise_int;
  wire [DATA_WIDTH - 1:0] qdr_q_fall_int;

  IDDR #(
    .DDR_CLK_EDGE ("SAME_EDGE_PIPELINED"),
    .INIT_Q1 (1'b0),
    .INIT_Q2 (1'b0),
    .SRTYPE ("SYNC")
  ) IDDR_qdrq [DATA_WIDTH - 1:0] (
    .C  (clk0),
    .CE (1'b1),
    .D  (qdr_q_iodelay),
    .R  (1'b0),
    .S  (1'b0),
    .Q1 (qdr_q_rise_int),
    .Q2 (qdr_q_fall_int)
  );

  assign qdr_q_rise = qdr_q_rise_int;
  assign qdr_q_fall = qdr_q_fall_int;

  /******************* SDR Inputs ********************
   * IODELAY for training
   */

endmodule
